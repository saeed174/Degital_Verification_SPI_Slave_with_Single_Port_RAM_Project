package shared_package;
    logic [2:0] next_mosi_shared  = 0;
    logic [10:0] old_MOSI_arr_shared = 0;
    int counter_shared  = 0;
endpackage