package shared_package;
    // logic [10:0] MOSI_arr_shared;
    // logic [2:0] next_mosi_shared  = 0;
    // logic [10:0] old_MOSI_arr_shared = 0;
    // int counter_shared  = 0;

    reg [2:0] cs_shared, ns_shared;
endpackage